`define COMMA_POSTV 10'b0101111100
`define COMMA_NEGTV 10'b1010000011