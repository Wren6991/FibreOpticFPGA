`timescale 1ns / 1ps

`define BIT_TIME 100

// Purpose: try all 2-symbol sequences
// and ensure that there are no runs of 5 or more bits.

module encode_8b10b_tb;

	// Inputs
	reg clk;
	reg rst;
	reg [7:0] d_in;
    reg nextword_enable;

	// Outputs
	wire [9:0] d_out;
	
	// Testvars for runlength-testing
	reg [19:0] d_out_history;
	reg t_fail;
	integer fail_count;
	integer i, j;

	// Instantiate the Unit Under Test (UUT)
	encode_8b10b uut (
		.clk(clk), 
		.rst(rst), 
		.d_in(d_in), 
		.d_out(d_out),
        .nextword_enable(nextword_enable),
		.idle(0)
	);

	always @ (posedge clk) begin
		d_out_history <= {d_out, d_out_history[19:10]};
		if (t_fail) begin
			fail_count <= fail_count + 1;
		end
	end

	// Generated with Python script lol
	always @ (*) begin
		/*
		// Check for run length
		casez (d_out_history)
			20'b11111???????????????: t_fail = 1;
			20'b?11111??????????????: t_fail = 1;
			20'b??11111?????????????: t_fail = 1;
			20'b???11111????????????: t_fail = 1;
			20'b????11111???????????: t_fail = 1;
			20'b?????11111??????????: t_fail = 1;
			20'b??????11111?????????: t_fail = 1;
			20'b???????11111????????: t_fail = 1;
			20'b????????11111???????: t_fail = 1;
			20'b?????????11111??????: t_fail = 1;
			20'b??????????11111?????: t_fail = 1;
			20'b???????????11111????: t_fail = 1;
			20'b????????????11111???: t_fail = 1;
			20'b?????????????11111??: t_fail = 1;
			20'b??????????????11111?: t_fail = 1;
			20'b???????????????11111: t_fail = 1;
			20'b00000???????????????: t_fail = 1;
			20'b?00000??????????????: t_fail = 1;
			20'b??00000?????????????: t_fail = 1;
			20'b???00000????????????: t_fail = 1;
			20'b????00000???????????: t_fail = 1;
			20'b?????00000??????????: t_fail = 1;
			20'b??????00000?????????: t_fail = 1;
			20'b???????00000????????: t_fail = 1;
			20'b????????00000???????: t_fail = 1;
			20'b?????????00000??????: t_fail = 1;
			20'b??????????00000?????: t_fail = 1;
			20'b???????????00000????: t_fail = 1;
			20'b????????????00000???: t_fail = 1;
			20'b?????????????00000??: t_fail = 1;
			20'b??????????????00000?: t_fail = 1;
			20'b???????????????00000: t_fail = 1;
			default: t_fail = 0;
		endcase*/
		
		// Check for comma sequence
		casez (d_out_history)
			20'b0101111100??????????: t_fail = 1;
			20'b?0101111100?????????: t_fail = 1;
			20'b??0101111100????????: t_fail = 1;
			20'b???0101111100???????: t_fail = 1;
			20'b????0101111100??????: t_fail = 1;
			20'b?????0101111100?????: t_fail = 1;
			20'b??????0101111100????: t_fail = 1;
			20'b???????0101111100???: t_fail = 1;
			20'b????????0101111100??: t_fail = 1;
			20'b?????????0101111100?: t_fail = 1;
			20'b??????????0101111100: t_fail = 1;
			20'b1010000011??????????: t_fail = 1;
			20'b?1010000011?????????: t_fail = 1;
			20'b??1010000011????????: t_fail = 1;
			20'b???1010000011???????: t_fail = 1;
			20'b????1010000011??????: t_fail = 1;
			20'b?????1010000011?????: t_fail = 1;
			20'b??????1010000011????: t_fail = 1;
			20'b???????1010000011???: t_fail = 1;
			20'b????????1010000011??: t_fail = 1;
			20'b?????????1010000011?: t_fail = 1;
			20'b??????????1010000011: t_fail = 1;
			default: t_fail = 0;
		endcase
	end


	always #(`BIT_TIME / 2) clk = ~clk;


	initial begin
		// Initialize Inputs
		clk = 1;
		rst = 1;
		d_in = 0;
		nextword_enable = 1;
		d_out_history = 0;
		fail_count = 0;

		// Wait 100 ns for global reset to finish
		#100;
		rst = 0;

		#(`BIT_TIME / 2)
		for (i = 0; i < 256; i = i + 1) begin
			for (j = 0; j < 256; j = j + 1) begin
				#`BIT_TIME
				d_in = i;
				#`BIT_TIME
				d_in = j;
				#`BIT_TIME
				d_in = i;
				#`BIT_TIME
				d_in = j;
			end
		end
        rst = 0;
        
		$finish;

	end
      
endmodule

