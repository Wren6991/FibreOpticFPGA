`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:50:54 05/21/2017 
// Design Name: 
// Module Name:    decode_8b10b 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

// Combinational circuit to decode 8b/10b non-control codewords
// Tables generated by python script lookup.py based on the 8b/10b Wikipedia article
module decode_8b10b(
    input [9:0] d_in,
    output reg [7:0] d_out
    );

always @(*) begin
    case (d_in[5:0])
        6'b100111: d_out[4:0] = 5'b00000;
        6'b011000: d_out[4:0] = 5'b00000;
        6'b011101: d_out[4:0] = 5'b00001;
        6'b100010: d_out[4:0] = 5'b00001;
        6'b101101: d_out[4:0] = 5'b00010;
        6'b010010: d_out[4:0] = 5'b00010;
        6'b110001: d_out[4:0] = 5'b00011;
        6'b110101: d_out[4:0] = 5'b00100;
        6'b001010: d_out[4:0] = 5'b00100;
        6'b101001: d_out[4:0] = 5'b00101;
        6'b011001: d_out[4:0] = 5'b00110;
        6'b111000: d_out[4:0] = 5'b00111;
        6'b000111: d_out[4:0] = 5'b00111;
        6'b111001: d_out[4:0] = 5'b01000;
        6'b000110: d_out[4:0] = 5'b01000;
        6'b100101: d_out[4:0] = 5'b01001;
        6'b010101: d_out[4:0] = 5'b01010;
        6'b110100: d_out[4:0] = 5'b01011;
        6'b001101: d_out[4:0] = 5'b01100;
        6'b101100: d_out[4:0] = 5'b01101;
        6'b011100: d_out[4:0] = 5'b01110;
        6'b010111: d_out[4:0] = 5'b01111;
        6'b101000: d_out[4:0] = 5'b01111;
        6'b011011: d_out[4:0] = 5'b10000;
        6'b100100: d_out[4:0] = 5'b10000;
        6'b100011: d_out[4:0] = 5'b10001;
        6'b010011: d_out[4:0] = 5'b10010;
        6'b110010: d_out[4:0] = 5'b10011;
        6'b001011: d_out[4:0] = 5'b10100;
        6'b101010: d_out[4:0] = 5'b10101;
        6'b011010: d_out[4:0] = 5'b10110;
        6'b111010: d_out[4:0] = 5'b10111;
        6'b000101: d_out[4:0] = 5'b10111;
        6'b110011: d_out[4:0] = 5'b11000;
        6'b001100: d_out[4:0] = 5'b11000;
        6'b100110: d_out[4:0] = 5'b11001;
        6'b010110: d_out[4:0] = 5'b11010;
        6'b110110: d_out[4:0] = 5'b11011;
        6'b001001: d_out[4:0] = 5'b11011;
        6'b001110: d_out[4:0] = 5'b11100;
        6'b101110: d_out[4:0] = 5'b11101;
        6'b010001: d_out[4:0] = 5'b11101;
        6'b011110: d_out[4:0] = 5'b11110;
        6'b100001: d_out[4:0] = 5'b11110;
        6'b101011: d_out[4:0] = 5'b11111;
        6'b010100: d_out[4:0] = 5'b11111;
        default: d_out[4:0] = 5'bxxxxx;
    endcase
    
    case (d_in[9:6])
        4'b1011: d_out[7:5] = 3'b000;
        4'b0100: d_out[7:5] = 3'b000;
        4'b1001: d_out[7:5] = 3'b001;
        4'b0101: d_out[7:5] = 3'b010;
        4'b1100: d_out[7:5] = 3'b011;
        4'b0011: d_out[7:5] = 3'b011;
        4'b1101: d_out[7:5] = 3'b100;
        4'b0010: d_out[7:5] = 3'b100;
        4'b1010: d_out[7:5] = 3'b101;
        4'b0110: d_out[7:5] = 3'b110;
        4'b1110: d_out[7:5] = 3'b111;
        4'b0001: d_out[7:5] = 3'b111;
        4'b0111: d_out[7:5] = 3'b111;
        4'b1000: d_out[7:5] = 3'b111;
        default: d_out[7:5] = 3'bxxx;
    endcase
end

endmodule
